`timescale 1ns / 1ps
`default_nettype none

module palette (
    input  wire       clk,
    input  wire [7:0] idx,
    output wire [8:0] pal_out
);

reg [8:0] data;

always @(posedge clk) begin case (idx)
    8'h00: data <= 9'b000000000;
    8'h01: data <= 9'b001000001;
    8'h02: data <= 9'b000000010;
    8'h03: data <= 9'b001000011;
    8'h04: data <= 9'b000000100;
    8'h05: data <= 9'b001000101;
    8'h06: data <= 9'b000000110;
    8'h07: data <= 9'b001000111;
    8'h08: data <= 9'b010000000;
    8'h09: data <= 9'b011000001;
    8'h0a: data <= 9'b010000010;
    8'h0b: data <= 9'b011000011;
    8'h0c: data <= 9'b010000100;
    8'h0d: data <= 9'b011000101;
    8'h0e: data <= 9'b010000110;
    8'h0f: data <= 9'b011000111;
    8'h10: data <= 9'b100000000;
    8'h11: data <= 9'b101000001;
    8'h12: data <= 9'b100000010;
    8'h13: data <= 9'b101000011;
    8'h14: data <= 9'b100000100;
    8'h15: data <= 9'b101000101;
    8'h16: data <= 9'b100000110;
    8'h17: data <= 9'b101000111;
    8'h18: data <= 9'b110000000;
    8'h19: data <= 9'b111000001;
    8'h1a: data <= 9'b110000010;
    8'h1b: data <= 9'b111000011;
    8'h1c: data <= 9'b110000100;
    8'h1d: data <= 9'b111000101;
    8'h1e: data <= 9'b110000110;
    8'h1f: data <= 9'b111000111;
    8'h20: data <= 9'b000001000;
    8'h21: data <= 9'b001001001;
    8'h22: data <= 9'b000001010;
    8'h23: data <= 9'b001001011;
    8'h24: data <= 9'b000001100;
    8'h25: data <= 9'b001001101;
    8'h26: data <= 9'b000001110;
    8'h27: data <= 9'b001001111;
    8'h28: data <= 9'b010001000;
    8'h29: data <= 9'b011001001;
    8'h2a: data <= 9'b010001010;
    8'h2b: data <= 9'b011001011;
    8'h2c: data <= 9'b010001100;
    8'h2d: data <= 9'b011001101;
    8'h2e: data <= 9'b010001110;
    8'h2f: data <= 9'b011001111;
    8'h30: data <= 9'b100001000;
    8'h31: data <= 9'b101001001;
    8'h32: data <= 9'b100001010;
    8'h33: data <= 9'b101001011;
    8'h34: data <= 9'b100001100;
    8'h35: data <= 9'b101001101;
    8'h36: data <= 9'b100001110;
    8'h37: data <= 9'b101001111;
    8'h38: data <= 9'b110001000;
    8'h39: data <= 9'b111001001;
    8'h3a: data <= 9'b110001010;
    8'h3b: data <= 9'b111001011;
    8'h3c: data <= 9'b110001100;
    8'h3d: data <= 9'b111001101;
    8'h3e: data <= 9'b110001110;
    8'h3f: data <= 9'b111001111;
    8'h40: data <= 9'b000010000;
    8'h41: data <= 9'b001010001;
    8'h42: data <= 9'b000010010;
    8'h43: data <= 9'b001010011;
    8'h44: data <= 9'b000010100;
    8'h45: data <= 9'b001010101;
    8'h46: data <= 9'b000010110;
    8'h47: data <= 9'b001010111;
    8'h48: data <= 9'b010010000;
    8'h49: data <= 9'b011010001;
    8'h4a: data <= 9'b010010010;
    8'h4b: data <= 9'b011010011;
    8'h4c: data <= 9'b010010100;
    8'h4d: data <= 9'b011010101;
    8'h4e: data <= 9'b010010110;
    8'h4f: data <= 9'b011010111;
    8'h50: data <= 9'b100010000;
    8'h51: data <= 9'b101010001;
    8'h52: data <= 9'b100010010;
    8'h53: data <= 9'b101010011;
    8'h54: data <= 9'b100010100;
    8'h55: data <= 9'b101010101;
    8'h56: data <= 9'b100010110;
    8'h57: data <= 9'b101010111;
    8'h58: data <= 9'b110010000;
    8'h59: data <= 9'b111010001;
    8'h5a: data <= 9'b110010010;
    8'h5b: data <= 9'b111010011;
    8'h5c: data <= 9'b110010100;
    8'h5d: data <= 9'b111010101;
    8'h5e: data <= 9'b110010110;
    8'h5f: data <= 9'b111010111;
    8'h60: data <= 9'b000011000;
    8'h61: data <= 9'b001011001;
    8'h62: data <= 9'b000011010;
    8'h63: data <= 9'b001011011;
    8'h64: data <= 9'b000011100;
    8'h65: data <= 9'b001011101;
    8'h66: data <= 9'b000011110;
    8'h67: data <= 9'b001011111;
    8'h68: data <= 9'b010011000;
    8'h69: data <= 9'b011011001;
    8'h6a: data <= 9'b010011010;
    8'h6b: data <= 9'b011011011;
    8'h6c: data <= 9'b010011100;
    8'h6d: data <= 9'b011011101;
    8'h6e: data <= 9'b010011110;
    8'h6f: data <= 9'b011011111;
    8'h70: data <= 9'b100011000;
    8'h71: data <= 9'b101011001;
    8'h72: data <= 9'b100011010;
    8'h73: data <= 9'b101011011;
    8'h74: data <= 9'b100011100;
    8'h75: data <= 9'b101011101;
    8'h76: data <= 9'b100011110;
    8'h77: data <= 9'b101011111;
    8'h78: data <= 9'b110011000;
    8'h79: data <= 9'b111011001;
    8'h7a: data <= 9'b110011010;
    8'h7b: data <= 9'b111011011;
    8'h7c: data <= 9'b110011100;
    8'h7d: data <= 9'b111011101;
    8'h7e: data <= 9'b110011110;
    8'h7f: data <= 9'b111011111;
    8'h80: data <= 9'b000100000;
    8'h81: data <= 9'b001100001;
    8'h82: data <= 9'b000100010;
    8'h83: data <= 9'b001100011;
    8'h84: data <= 9'b000100100;
    8'h85: data <= 9'b001100101;
    8'h86: data <= 9'b000100110;
    8'h87: data <= 9'b001100111;
    8'h88: data <= 9'b010100000;
    8'h89: data <= 9'b011100001;
    8'h8a: data <= 9'b010100010;
    8'h8b: data <= 9'b011100011;
    8'h8c: data <= 9'b010100100;
    8'h8d: data <= 9'b011100101;
    8'h8e: data <= 9'b010100110;
    8'h8f: data <= 9'b011100111;
    8'h90: data <= 9'b100100000;
    8'h91: data <= 9'b101100001;
    8'h92: data <= 9'b100100010;
    8'h93: data <= 9'b101100011;
    8'h94: data <= 9'b100100100;
    8'h95: data <= 9'b101100101;
    8'h96: data <= 9'b100100110;
    8'h97: data <= 9'b101100111;
    8'h98: data <= 9'b110100000;
    8'h99: data <= 9'b111100001;
    8'h9a: data <= 9'b110100010;
    8'h9b: data <= 9'b111100011;
    8'h9c: data <= 9'b110100100;
    8'h9d: data <= 9'b111100101;
    8'h9e: data <= 9'b110100110;
    8'h9f: data <= 9'b111100111;
    8'ha0: data <= 9'b000101000;
    8'ha1: data <= 9'b001101001;
    8'ha2: data <= 9'b000101010;
    8'ha3: data <= 9'b001101011;
    8'ha4: data <= 9'b000101100;
    8'ha5: data <= 9'b001101101;
    8'ha6: data <= 9'b000101110;
    8'ha7: data <= 9'b001101111;
    8'ha8: data <= 9'b010101000;
    8'ha9: data <= 9'b011101001;
    8'haa: data <= 9'b010101010;
    8'hab: data <= 9'b011101011;
    8'hac: data <= 9'b010101100;
    8'had: data <= 9'b011101101;
    8'hae: data <= 9'b010101110;
    8'haf: data <= 9'b011101111;
    8'hb0: data <= 9'b100101000;
    8'hb1: data <= 9'b101101001;
    8'hb2: data <= 9'b100101010;
    8'hb3: data <= 9'b101101011;
    8'hb4: data <= 9'b100101100;
    8'hb5: data <= 9'b101101101;
    8'hb6: data <= 9'b100101110;
    8'hb7: data <= 9'b101101111;
    8'hb8: data <= 9'b110101000;
    8'hb9: data <= 9'b111101001;
    8'hba: data <= 9'b110101010;
    8'hbb: data <= 9'b111101011;
    8'hbc: data <= 9'b110101100;
    8'hbd: data <= 9'b111101101;
    8'hbe: data <= 9'b110101110;
    8'hbf: data <= 9'b111101111;
    8'hc0: data <= 9'b000110000;
    8'hc1: data <= 9'b001110001;
    8'hc2: data <= 9'b000110010;
    8'hc3: data <= 9'b001110011;
    8'hc4: data <= 9'b000110100;
    8'hc5: data <= 9'b001110101;
    8'hc6: data <= 9'b000110110;
    8'hc7: data <= 9'b001110111;
    8'hc8: data <= 9'b010110000;
    8'hc9: data <= 9'b011110001;
    8'hca: data <= 9'b010110010;
    8'hcb: data <= 9'b011110011;
    8'hcc: data <= 9'b010110100;
    8'hcd: data <= 9'b011110101;
    8'hce: data <= 9'b010110110;
    8'hcf: data <= 9'b011110111;
    8'hd0: data <= 9'b100110000;
    8'hd1: data <= 9'b101110001;
    8'hd2: data <= 9'b100110010;
    8'hd3: data <= 9'b101110011;
    8'hd4: data <= 9'b100110100;
    8'hd5: data <= 9'b101110101;
    8'hd6: data <= 9'b100110110;
    8'hd7: data <= 9'b101110111;
    8'hd8: data <= 9'b110110000;
    8'hd9: data <= 9'b111110001;
    8'hda: data <= 9'b110110010;
    8'hdb: data <= 9'b111110011;
    8'hdc: data <= 9'b110110100;
    8'hdd: data <= 9'b111110101;
    8'hde: data <= 9'b110110110;
    8'hdf: data <= 9'b111110111;
    8'he0: data <= 9'b000111000;
    8'he1: data <= 9'b001111001;
    8'he2: data <= 9'b000111010;
    8'he3: data <= 9'b001111011;
    8'he4: data <= 9'b000111100;
    8'he5: data <= 9'b001111101;
    8'he6: data <= 9'b000111110;
    8'he7: data <= 9'b001111111;
    8'he8: data <= 9'b010111000;
    8'he9: data <= 9'b011111001;
    8'hea: data <= 9'b010111010;
    8'heb: data <= 9'b011111011;
    8'hec: data <= 9'b010111100;
    8'hed: data <= 9'b011111101;
    8'hee: data <= 9'b010111110;
    8'hef: data <= 9'b011111111;
    8'hf0: data <= 9'b100111000;
    8'hf1: data <= 9'b101111001;
    8'hf2: data <= 9'b100111010;
    8'hf3: data <= 9'b101111011;
    8'hf4: data <= 9'b100111100;
    8'hf5: data <= 9'b101111101;
    8'hf6: data <= 9'b100111110;
    8'hf7: data <= 9'b101111111;
    8'hf8: data <= 9'b110111000;
    8'hf9: data <= 9'b111111001;
    8'hfa: data <= 9'b110111010;
    8'hfb: data <= 9'b111111011;
    8'hfc: data <= 9'b110111100;
    8'hfd: data <= 9'b111111101;
    8'hfe: data <= 9'b110111110;
    8'hff: data <= 9'b111111111;
endcase end
    
assign pal_out = data;

endmodule

`default_nettype wire