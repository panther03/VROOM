`define KONATA_ENABLE
//`define DEBUG_ENABLE